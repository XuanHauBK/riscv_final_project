//-----------------------------------------------------------------------------
//    Copyright (C) 2016 by Dolphin Technology
//    All right reserved.
//    
//    Copyright Notification
//    No part may be reproduced except as authorized by written permission.
//    
//    File: ../hdl/rb_derivative_reg.sv
//    Project: dti_uart
//    Author: hautx0
//    Created: Sep 23rd 2024
//    Description:
//       Derivative Registers
//    
//    History:
//    Date ------------ By ------------ Change Description
//------------------------------------------------------------------------------
module rb_derivative_reg ( 
// Field Signals
// Derivative Signals
// End
);

//-------------------------------------------------------------------------
// Assignments
//-------------------------------------------------------------------------

endmodule